*
.SUBCKT LT1008 3 2 7 4 6 1 8
* USE C=30 PF IN MAIN CIRCUIT (CA TO CB).
* INPUT
RC1 7 80 8842
RC2 7 90 8842
Q1 80 2 10 QM1
Q2 90 3 11 QM2
DDM1 2 3 DM2
DDM2 3 2 DM2
C1 80 90 8.66e-12
RE1 10 12 224.6
RE2 11 12 224.6
IEE 12 4 6e-6
RE 12 0 33330000
CE 12 0 1.579E-12
* INTERMEDIATE
GCM 0 8 12 0 2.841E-11
GA 8 0 80 90 1.131E-04
R2 8 0 100000
* EXTERNAL COMP CAP USED FOR C2 (SEE NOTE ABOVE).
GB 1 0 8 0 196
* OUTPUT
RO1 1 6 100
RO2 1 0 900
RC 17 0 6.802e-5
GC 0 17 6 0 14700
D1 1 17 DM1
D2 17 1 DM1
D3 6 13 DM2
D4 14 6 DM2
VC 7 13 1.774
VE 14 4 1.774
IP 7 4 0.000374
DSUB 4 7 DM2
.MODEL QM1 NPN(IS=8e-16 BF=66670)
.MODEL QM2 NPN(IS=8.009E-16 BF=200000)
.MODEL DM1 D(IS=4.276E-12)
.MODEL DM2 D(IS=8e-16)
.ENDS LT1008
XU1 0 4 3 7 6 2 1 LT1008
V1 0 7 15
V2 3 0 15
V3 5 0 SINE(0 0.1 1k)
R2 4 5 2k
R1 6 4 7k
C1 0 0 30p
* INSTRUCTIONS: Check that your 1 kHz sinusoidal input voltage amplitude is below 100mV and the output voltage is also sinusoidal (not slew rate limited). Measure the gain.
* SIMULATION NOTES: For the purposes of simulation, set the amplitude of the input signal to exactly 100mV. The simulation time should be 2 milliseconds
* CODE: 111A
.control
tran 5u 2m
run
print v(4) v(5)
.endc