*** Ammeter Connected to first position, Q3 Q4 Base Grounded via Jumper ***
.subckt CA3083 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
Q3 1 16 15 QM1
Q1 2 3 4 QM1
Q2 7 6 8 QM1
Q4 9 10 11 QM1
Q5 14 13 12 QM1
.MODEL QM1 NPN(IS=8e-16 BF=66670)
.ends CA3083
XU1 7 8 11 9 0 9 3 4 3 3 4 0 0 0 10 9 CA3083
RB 2 3 1k
C1 0 0 30p
RC1 5 7 1k
RC2 6 8 1k
R4a 0 0 4k
R4b 0 0 4k
R3a 0 0 4k
R3a 0 0 4k
R2 0 0 4k
R7 0 0 4k
R8 0 0 4k
R9 0 0 4k
V1 1 0 dc 1
V2 0 4 dc 1
RAmmeter1 1 2 1m
RJumper1 1 5 1m
RJumper2 1 6 1m
RJumper3 0 0 1m
RJumper4 10 0 10m
RJumper5 11 0 1m
XU2 13 12 0 0 14 LM741
.MODEL QM1 NPN(IS=8e-16 BF=66670)
* INSTRUCTIONS: Creative mode allows you to construct, simulate and implement a circuit in any way within the constraints of the hardware. You have been provided with every node necessary for constructing the circuit. Joining nodes will produce an error.
* IMPLEMENTATION NOTES: When this lab is opened, the relay controlling the power supply (Power - Port 1 Line 3 - ON) will switch ON. Once your circuit has been constructed, it will be checked against a set of possible valid implementations. If your circuit matches, it will be implemented on the hardware
* DIGOUTPUT0_PRE = 0 1 1 0 0 0 0 0
* DIGOUTPUT1_PRE = 0 0 0 1 0 0 0 0
* DIGOUTPUT0_POST = 1 0 0 0 0 0 0 0
* DIGOUTPUT1_POST = 0 0 0 1 0 0 0 0
* AOUTPUT0_PRE = 0.0
* AOUTPUT1_PRE = 0.0
* AOUTPUT0_POST = 0.0 
* AOUTPUT1_POST = 0.0
*** Ammeter Connected to second position, Q3 Q4 Base Grounded via Jumper ***
XU1 7 8 10 9 0 3 3 4 9 3 4 0 0 0 9 0 CA3083
RB 2 3 1k
C1 0 0 30p
RC1 5 7 1k
RC2 6 8 1k
R4a 0 0 4k
R4b 0 0 4k
R3a 0 0 4k
R3a 0 0 4k
R2 0 0 4k
R7 0 0 4k
R8 0 0 4k
R9 0 0 4k
V1 1 0 dc 1
V2 0 4 dc 1
RAmmeter1 1 2 1m
RJumper1 1 5 1m
RJumper2 1 6 1m
RJumper3 0 0 1m
XU2 11 10 1 4 12 LM741
.MODEL QM1 NPN(IS=8e-16 BF=66670)
* INSTRUCTIONS: Creative mode allows you to construct, simulate and implement a circuit in any way within the constraints of the hardware. You have been provided with every node necessary for constructing the circuit. Joining nodes will produce an error.
* IMPLEMENTATION NOTES: When this lab is opened, the relay controlling the power supply (Power - Port 1 Line 3 - ON) will switch ON. Once your circuit has been constructed, it will be checked against a set of possible valid implementations. If your circuit matches, it will be implemented on the hardware
* DIGOUTPUT0_PRE = 0 1 1 0 0 0 0 0
* DIGOUTPUT1_PRE = 0 0 0 1 0 0 0 0
* DIGOUTPUT0_POST = 1 0 0 0 0 0 0 0
* DIGOUTPUT1_POST = 0 0 0 1 0 0 0 0
* AOUTPUT0_PRE = 0.0
* AOUTPUT1_PRE = 0.0
* AOUTPUT0_POST = 0.0 
* AOUTPUT1_POST = 0.0
*** Ammeter Connected to third position, Q3 Q4 Base Grounded via Jumper ***
XU1 7 8 0 9 0 3 3 4 9 3 4 0 0 0 9 0 CA3083
RB 2 3 1k
C1 0 0 30p
RC1 5 7 1k
RC2 6 8 1k
R4a 0 0 4k
R4b 0 0 4k
R3a 0 0 4k
R3a 0 0 4k
R2 0 0 4k
R7 0 0 4k
R8 0 0 4k
R9 0 0 4k
V1 1 0 dc 1
V2 0 4 dc 1
RAmmeter1 1 2 1m
RJumper1 1 5 1m
RJumper2 1 6 1m
RJumper3 0 0 1m
XU2 11 10 1 4 12 LM741
.MODEL QM1 NPN(IS=8e-16 BF=66670)
* INSTRUCTIONS: Creative mode allows you to construct, simulate and implement a circuit in any way within the constraints of the hardware. You have been provided with every node necessary for constructing the circuit. Joining nodes will produce an error.
* IMPLEMENTATION NOTES: When this lab is opened, the relay controlling the power supply (Power - Port 1 Line 3 - ON) will switch ON. Once your circuit has been constructed, it will be checked against a set of possible valid implementations. If your circuit matches, it will be implemented on the hardware
* DIGOUTPUT0_PRE = 0 1 1 0 0 0 0 0
* DIGOUTPUT1_PRE = 0 0 0 1 0 0 0 0
* DIGOUTPUT0_POST = 1 0 0 0 0 0 0 0
* DIGOUTPUT1_POST = 0 0 0 1 0 0 0 0
* AOUTPUT0_PRE = 0.0
* AOUTPUT1_PRE = 0.0
* AOUTPUT0_POST = 0.0 
* AOUTPUT1_POST = 0.0
*** No Ammeter, Signal Generator 1kHz at Input ***
XU1 7 8 0 9 0 3 3 4 9 3 4 0 0 0 9 0 CA3083
RB 2 3 1k
C1 0 0 30p
RC1 5 7 1k
RC2 6 8 1k
R4a 0 0 4k
R4b 0 0 4k
R3a 0 0 4k
R3a 0 0 4k
R2 0 0 4k
R7 0 0 4k
R8 0 0 4k
R9 0 0 4k
V1 1 0 dc 1
V2 0 4 dc 1
V3 9 0 SINE(0 4m 1k)
RAmmeter1 0 0 1m
RJumper1 1 2 1m
RJumper2 1 5 1m
RJumper3 1 6 1m
XU2 11 10 1 4 12 LM741
.MODEL QM1 NPN(IS=8e-16 BF=66670)
* INSTRUCTIONS: Creative mode allows you to construct, simulate and implement a circuit in any way within the constraints of the hardware. You have been provided with every node necessary for constructing the circuit. Joining nodes will produce an error.
* IMPLEMENTATION NOTES: When this lab is opened, the relay controlling the power supply (Power - Port 1 Line 3 - ON) will switch ON. Once your circuit has been constructed, it will be checked against a set of possible valid implementations. If your circuit matches, it will be implemented on the hardware
* DIGOUTPUT0_PRE = 0 1 1 0 0 0 0 0
* DIGOUTPUT1_PRE = 0 0 0 1 0 0 0 0
* DIGOUTPUT0_POST = 1 0 0 0 0 0 0 0
* DIGOUTPUT1_POST = 0 0 0 1 0 0 0 0
* AOUTPUT0_PRE = 0.0
* AOUTPUT1_PRE = 0.0
* AOUTPUT0_POST = 0.0 
* AOUTPUT1_POST = 0.0
*** No Ammeter, Signal Generator 1kHz at Input and Capacitor ***
XU1 7 8 0 9 0 3 3 4 9 3 4 0 0 0 9 0 CA3083
RB 2 3 1k
C1 7 8 30p
RC1 5 7 1k
RC2 6 8 1k
R4a 0 0 4k
R4b 0 0 4k
R3a 0 0 4k
R3a 0 0 4k
R2 0 0 4k
R7 0 0 4k
R8 0 0 4k
R9 0 0 4k
V1 1 0 dc 1
V2 0 4 dc 1
V3 9 0 SINE(0 4m 1k)
RAmmeter1 0 0 1m
RJumper1 1 2 1m
RJumper2 1 5 1m
RJumper3 1 6 1m
XU2 11 10 1 4 12 LM741
.MODEL QM1 NPN(IS=8e-16 BF=66670)
* INSTRUCTIONS: Creative mode allows you to construct, simulate and implement a circuit in any way within the constraints of the hardware. You have been provided with every node necessary for constructing the circuit. Joining nodes will produce an error.
* IMPLEMENTATION NOTES: When this lab is opened, the relay controlling the power supply (Power - Port 1 Line 3 - ON) will switch ON. Once your circuit has been constructed, it will be checked against a set of possible valid implementations. If your circuit matches, it will be implemented on the hardware
* DIGOUTPUT0_PRE = 0 1 1 0 0 0 0 0
* DIGOUTPUT1_PRE = 0 0 0 1 0 0 0 0
* DIGOUTPUT0_POST = 1 0 0 0 0 0 0 0
* DIGOUTPUT1_POST = 0 0 0 1 0 0 0 0
* AOUTPUT0_PRE = 0.0
* AOUTPUT1_PRE = 0.0
* AOUTPUT0_POST = 0.0 
* AOUTPUT1_POST = 0.0
*** No Ammeter, Signal Generator 1kHz at Input and Capacitor ***
XU1 7 8 0 9 0 3 3 4 9 3 4 0 0 0 9 0 CA3083
RB 2 3 1k
C1 7 8 30p
RC1 5 7 1k
RC2 6 8 1k
R4a 0 0 4k
R4b 0 0 4k
R3a 0 0 4k
R3a 0 0 4k
R2 0 0 4k
R7 0 0 4k
R8 0 0 4k
R9 0 0 4k
V1 1 0 dc 1
V2 0 4 dc 1
V3 9 0 SINE(0 4m 1k)
RAmmeter1 0 0 1m
RJumper1 1 2 1m
RJumper2 1 5 1m
RJumper3 1 6 1m
XU2 11 10 1 4 12 LM741
.MODEL QM1 NPN(IS=8e-16 BF=66670)
* INSTRUCTIONS: Creative mode allows you to construct, simulate and implement a circuit in any way within the constraints of the hardware. You have been provided with every node necessary for constructing the circuit. Joining nodes will produce an error.
* IMPLEMENTATION NOTES: When this lab is opened, the relay controlling the power supply (Power - Port 1 Line 3 - ON) will switch ON. Once your circuit has been constructed, it will be checked against a set of possible valid implementations. If your circuit matches, it will be implemented on the hardware
* DIGOUTPUT0_PRE = 0 1 1 0 0 0 0 0
* DIGOUTPUT1_PRE = 0 0 0 1 0 0 0 0
* DIGOUTPUT0_POST = 1 0 0 0 0 0 0 0
* DIGOUTPUT1_POST = 0 0 0 1 0 0 0 0
* AOUTPUT0_PRE = 0.0
* AOUTPUT1_PRE = 0.0
* AOUTPUT0_POST = 0.0 
* AOUTPUT1_POST = 0.0