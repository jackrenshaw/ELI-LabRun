* /Users/jackrenshaw/dev/ELI/labs/Amplifier with Feedback/Part A: Differential Amplifier/Draft1.asc
V1 N001 0 15V
Q1 N007 N007 N010 0 NPN
R1 N001 N007 1k
Q2 N004 N006 N008 0 NPN
Q3 N002 N005 N008 0 NPN
Q4 N008 N007 N010 0 NPN
R2 N001 N002 1k
R3 N001 N004 1k
R4 N009 0 1k
V2 N005 0 SINE(0 1 1k)
C1 N004 N002 100p
R5 N004 0 1k
R6 N003 N002 1k
R7 N003 N009 1k
V3 0 N010 15V
.model NPN NPN
.model PNP PNP
.tran 50u 500m
.control
tran 50u 500m
run
print v(N002)
.endc