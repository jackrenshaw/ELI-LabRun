*
.SUBCKT LM348N  1 2 3 4 5 6 7 8 9 10 11 12 13 14
* Dummy subcircuit, can someone please develop?!
.ENDS LM348N
.MODEL d1 D(IS=18.8n RS=0 BV=400 IBV=5u CJO=30 M=0.333 N=2)
XA 1 999 999 4 0 7 7 8 0 10 11 0 13 14 LM348N
RVariable1 4 5 10k
RVariable2 5 11 10k
C1 6 7 10p
Rx11 7 10 1k
Rx12 7 10 1k
Rx13 7 10 1k
Rx14 7 10 1k
Rx15 7 10 1k
Rx16 7 10 1k
R21 10 8 1k
R31 2 6 1k
R32 2 6 1k
V1 4 0 15
V2 0 11 15
V3 999 0 0
* INSTRUCTIONS: Creative mode allows you to construct, simulate and implement a circuit in any way within the constraints of the hardware. You have been provided with every node necessary for constructing the circuit. Joining nodes will produce an error.
* IMPLEMENTATION NOTES: When this lab is opened, the relay controlling the power supply (Power - Port 1 Line 3 - ON) will switch ON. Once your circuit has been constructed, it will be checked against a set of possible valid implementations. If your circuit matches, it will be implemented on the hardware
* DIGOUTPUT0_PRE = 0 0 0 0 0 0 0 0
* DIGOUTPUT1_PRE = 0 0 0 0 0 0 0 0
* AOUTPUT0_PRE = 0.0
* AOUTPUT1_PRE = 0.0
.control
tran 20u 1m
run
print v(6)
dc V1 15 15 0.1
dc V2 15 15 0.1
run
print v(11) v(4) v(5)
.endc