*
.subckt lm741 Pin1_IN_$$PLUS$ Pin2_IN_$$MINUS$
+ Pin3_V_$$PLUS$ Pin4_V_$$MINUS$ Pin5_OUT
RU2$U4$R1 Pin4_V_$$MINUS$ U2$U4$OUT 144.0
RU2$U4$R2 U2$U4$OUT Pin3_V_$$PLUS$ 144.0
DU2$U4$D6 U2$U4$DRIVE_OUT U2$U4$V1_PIN_1 DG1 temp=27
.model DG1 D IS=1.0E-12
RU2$U4$R36 U2$U4$DRIVE_OUT Pin4_V_$$MINUS$ 2000000.0
RU2$U4$R38 Pin3_V_$$PLUS$ U2$U4$DRIVE_OUT 2000000.0
DU2$U4$D4 Pin3_V_$$PLUS$ U2$U4$D2_PIN_2 DG2
.model DG2 D
DU2$U4$D5 Pin4_V_$$MINUS$ U2$U4$D3_PIN_2 DG3
.model DG3 D BV=50.0
DU2$U4$D3 Pin3_V_$$PLUS$ U2$U4$D3_PIN_2 DG4
.model DG4 D
DU2$U4$D1 U2$U4$D1_PIN_1 U2$U4$DRIVE_OUT DG5 temp=27
.model DG5 D IS=1.0E-12
DU2$U4$D2 Pin4_V_$$MINUS$ U2$U4$D2_PIN_2 DG6
.model DG6 D BV=50.0
GU2$U4$B2$controlledSource U2$U4$D2_PIN_2 Pin4_V_$$MINUS$
+ VALUE={V(U2$U4$DRIVE_OUT, U2$U4$OUT) / (2.0 * 72.0)}
GU2$U4$G2$3 U2$U4$OUT Pin4_V_$$MINUS$ VALUE={-1.0 / (2.0 *
+ 72.0) * V(U2$U4$DRIVE_OUT, Pin4_V_$$MINUS$)}
VU2$U4$V2$1 U2$U4$OUT U2$U4$D1_PIN_1 1.3426910213823116
GU2$U4$B1$controlledSource U2$U4$D3_PIN_2 Pin4_V_$$MINUS$
+ VALUE={V(U2$U4$OUT, U2$U4$DRIVE_OUT) / (2.0 * 72.0)}
LU2$U4$L1$inductor U2$U4$L1$currentProbe$_PIN1 U2$U4$OUT
+ 5.0E-7 IC=0.0
VU2$U4$L1$resistor U2$U4$L1$currentProbe$_PIN2 Pin5_OUT
+ 0.0
VU2$U4$L1$currentProbe U2$U4$L1$currentProbe$_PIN1
+ U2$U4$L1$currentProbe$_PIN2 0
VU2$U4$V1$1 U2$U4$V1_PIN_1 U2$U4$OUT 1.3426910213823116
GU2$U4$B6$controlledSource Pin4_V_$$MINUS$ U2$U4$DRIVE_OUT
+ VALUE={(V(Pin3_V_$$PLUS$, Pin4_V_$$MINUS$) / 2.0 +
+ V(U2$U9$Pin_2_OUT)) / (2.0 * 1000000.0)}
GU2$U4$G1$3 Pin3_V_$$PLUS$ U2$U4$OUT VALUE={-1.0 / (2.0 *
+ 72.0) * V(Pin3_V_$$PLUS$, U2$U4$DRIVE_OUT)}
GU2$U4$B5$controlledSource U2$U4$DRIVE_OUT Pin3_V_$$PLUS$
+ VALUE={(V(Pin3_V_$$PLUS$, Pin4_V_$$MINUS$) / 2.0 -
+ V(U2$U9$Pin_2_OUT)) / (2.0 * 1000000.0)}
RU2$U2$R39 U2$U2$L1_PIN_1 0 10000.0
RU2$U2$U2$R40 U2$U2$U2$R39_PIN_1 U2$U2$U2$Q2_PIN_3
+ 0.8109886183790636
RU2$U2$U2$R1 U2$U5$Pin_2_IN_$$MINUS$ Pin3_V_$$PLUS$
+ 31.830988618379063
RU2$U2$U2$R2 U2$U5$Pin_1_IN_$$PLUS$ Pin3_V_$$PLUS$
+ 31.830988618379063
QU2$U2$U2$Q1 U2$U5$Pin_2_IN_$$MINUS$
+ U2$U2$U2$Pin_1_IN_$$PLUS$ U2$U2$U2$R39_PIN_2 QG7 OFF
.model QG7 NPN BF=15151.515151515152
QU2$U2$U2$Q2 U2$U5$Pin_1_IN_$$PLUS$ Pin2_IN_$$MINUS$
+ U2$U2$U2$Q2_PIN_3 QG8 OFF
.model QG8 NPN BF=15151.515151515152
RU2$U2$U2$R39 U2$U2$U2$R39_PIN_1 U2$U2$U2$R39_PIN_2
+ 0.8109886183790636
IU2$U2$U2$I1$1 U2$U2$U2$R39_PIN_1 Pin4_V_$$MINUS$
+ 0.0016666666666666668
GU2$U2$I4$controlledSource 0 U2$U2$F_VCM_CMRR
+ VALUE={((V(Pin1_IN_$$PLUS$) + V(Pin2_IN_$$MINUS$)) / 2.0 -
+ (V(Pin3_V_$$PLUS$) + V(Pin4_V_$$MINUS$)) / 2.0) / 10000.0
+ / 30000.0}
LU2$U2$L1$inductor U2$U2$L1$currentProbe$_PIN1
+ U2$U2$L1_PIN_1 5.305164769729845 IC=0.0
VU2$U2$L1$resistor U2$U2$L1$currentProbe$_PIN2
+ U2$U2$F_VCM_CMRR 0.0
VU2$U2$L1$currentProbe U2$U2$L1$currentProbe$_PIN1
+ U2$U2$L1$currentProbe$_PIN2 0
EU2$U2$V11$controlledSource U2$U2$U2$Pin_1_IN_$$PLUS$
+ Pin1_IN_$$PLUS$ VALUE={0.0 + V(U2$U2$F_VCM_CMRR)}
IU2$U2$I5$1 Pin1_IN_$$PLUS$ Pin2_IN_$$MINUS$ 0.0
CU2$U2$C8$1 Pin1_IN_$$PLUS$ U2$U2$C8$2$_PIN1 1.5E-12
+ IC=0.0
VU2$U2$C8$2 U2$U2$C8$2$_PIN1 Pin2_IN_$$MINUS$ 0.0
CU2$U2$C9$1 U2$U5$Pin_2_IN_$$MINUS$ U2$U2$C9$2$_PIN1
+ 2.0798668885191352E-10 IC=0.0
VU2$U2$C9$2 U2$U2$C9$2$_PIN1 U2$U5$Pin_1_IN_$$PLUS$ 0.0
RU2$U6$R1 0 U2$U7$Pin_1_IN 1000000.0
GU2$U6$G1$3 0 U2$U7$Pin_1_IN VALUE={1.0 / 1000000.0 *
+ V(U2$U5$Pin_5_OUT, 0)}
CU2$U6$C1$1 0 U2$U6$C1$2$_PIN1 1.3240843851239214E-14
+ IC=0.0
VU2$U6$C1$2 U2$U6$C1$2$_PIN1 U2$U7$Pin_1_IN 0.0
RU2$U8$R1 0 U2$U9$Pin_1_IN 1000000.0
GU2$U8$G1$3 0 U2$U9$Pin_1_IN VALUE={1.0 / 1000000.0 *
+ V(U2$U7$Pin_2_OUT, 0)}
CU2$U8$C1$1 0 U2$U8$C1$2$_PIN1 1.3240843851239214E-14
+ IC=0.0
VU2$U8$C1$2 U2$U8$C1$2$_PIN1 U2$U9$Pin_1_IN 0.0
RU2$U9$R1 0 U2$U9$Pin_2_OUT 1000000.0
GU2$U9$G1$3 0 U2$U9$Pin_2_OUT VALUE={1.0 / 1000000.0 *
+ V(U2$U9$Pin_1_IN, 0)}
CU2$U9$C1$1 0 U2$U9$C1$2$_PIN1 1.3240843851239214E-14
+ IC=0.0
VU2$U9$C1$2 U2$U9$C1$2$_PIN1 U2$U9$Pin_2_OUT 0.0
RU2$U7$R1 0 U2$U7$Pin_2_OUT 1000000.0
GU2$U7$G1$3 0 U2$U7$Pin_2_OUT VALUE={1.0 / 1000000.0 *
+ V(U2$U7$Pin_1_IN, 0)}
CU2$U7$C1$1 0 U2$U7$C1$2$_PIN1 1.3240843851239214E-14
+ IC=0.0
VU2$U7$C1$2 U2$U7$C1$2$_PIN1 U2$U7$Pin_2_OUT 0.0
DU2$U5$D9 U2$U5$Pin_5_OUT U2$U5$V10_PIN_2 DG9 temp=27
.model DG9 D IS=1.0E-12
RU2$U5$R36 0 U2$U5$Pin_5_OUT 477464.82927568594
DU2$U5$D10 U2$U5$D10_PIN_1 U2$U5$Pin_5_OUT DG10 temp=27
.model DG10 D IS=1.0E-12
EU2$U5$V8$controlledSource U2$U5$V10_PIN_1 0
+ VALUE={V(Pin3_V_$$PLUS$, Pin4_V_$$MINUS$) / 2.0}
EU2$U5$B3$controlledSource 0 U2$U5$V9_PIN_2
+ VALUE={V(Pin3_V_$$PLUS$, Pin4_V_$$MINUS$) / 2.0}
CU2$U5$C5$1 0 U2$U5$C5$2$_PIN1 3.3333333333333334E-9
+ IC=0.0
VU2$U5$C5$2 U2$U5$C5$2$_PIN1 U2$U5$Pin_5_OUT 0.0
GU2$U5$G7$3 0 U2$U5$Pin_5_OUT VALUE={15000.0 /
+ 477464.82927568594 * V(U2$U5$Pin_1_IN_$$PLUS$,
+ U2$U5$Pin_2_IN_$$MINUS$)}
VU2$U5$V9$1 U2$U5$D10_PIN_1 U2$U5$V9_PIN_2
+ 1.5489012642594155
VU2$U5$V10$1 U2$U5$V10_PIN_1 U2$U5$V10_PIN_2
+ 1.5489012642594155
.ends lm741
* This is the potentiometer
*      _____
*  1--|_____|--2
*        |
*        3
*
.MODEL d1 D(IS=18.8n RS=0 BV=400 IBV=5u CJO=30 M=0.333 N=2)
* XA 5 2 4 11 1 LM741
XB 0 6 4 11 6 LM741
XC 10 9 4 11 8 LM741
* XD 12 13 4 11 14 LM741
RVariable1 4 5 100k
RVariable2 5 11 100k
Rx11 6 10 1k
Rx12 6 10 1k
Rx13 6 10 1k
Rx14 6 10 1k
Rx15 6 10 1k
Rx16 6 10 1k
R21 10 8 1k
V1 4 0 15
V2 0 11 15
V3 999 999 0
C 6 7 10p
R41 8 2 1k
R32 2 6 1k
R31 999 999 1k
* INSTRUCTIONS: Creative mode allows you to construct, simulate and implement a circuit in any way within the constraints of the hardware. You have been provided with every node necessary for constructing the circuit. Joining nodes will produce an error.
* IMPLEMENTATION NOTES: When this lab is opened, the relay controlling the power supply (Power - Port 1 Line 3 - ON) will switch ON. Once your circuit has been constructed, it will be checked against a set of possible valid implementations. If your circuit matches, it will be implemented on the hardware
* DIGOUTPUT0_PRE = 0 0 0 0 0 0 0 0
* DIGOUTPUT1_PRE = 0 0 0 0 0 0 0 0
* DIGOUTPUT0_POST = 0 0 0 0 0 0 0 0
* DIGOUTPUT1_POST = 0 0 0 0 0 0 0 0
* AOUTPUT0_PRE = 0.0
* AOUTPUT1_PRE = 0.0
* AOUTPUT0_POST = 0.0 
* AOUTPUT1_POST = 0.0
* AOUTPUT0_DEVICE = RVariable1
* AOUTPUT0_MINV = 0.0
* AOUTPUT0_MAXV = 5.0
* AOUTPUT1_DEVICE = RVariable1
* AOUTPUT1_MINV = 0.0
* AOUTPUT1_MAXV = 5.0
.control
tran 20u 20m
run
print v(7) v(10)
dc V1 15 15 0.1
dc V2 15 15 0.1
run
print v(1) v(2) v(3) v(4) v(5) v(6) v(7) V(8) v(9) v(10) v(11) v(12) v(13) v(14) v(15)
.endc