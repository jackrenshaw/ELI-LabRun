*
.SUBCKT LT1008 3 2 7 4 6 1 8
* USE C=30 PF IN MAIN CIRCUIT (CA TO CB).
* INPUT
RC1 7 80 8842
RC2 7 90 8842
Q1 80 2 10 QM1
Q2 90 3 11 QM2
DDM1 2 3 DM2
DDM2 3 2 DM2
C1 80 90 8.66e-12
RE1 10 12 224.6
RE2 11 12 224.6
IEE 12 4 6e-6
RE 12 0 33330000
CE 12 0 1.579E-12
* INTERMEDIATE
GCM 0 8 12 0 2.841E-11
GA 8 0 80 90 1.131E-04
R2 8 0 100000
* EXTERNAL COMP CAP USED FOR C2 (SEE NOTE ABOVE).
GB 1 0 8 0 196
* OUTPUT
RO1 1 6 100
RO2 1 0 900
RC 17 0 6.802e-5
GC 0 17 6 0 14700
D1 1 17 DM1
D2 17 1 DM1
D3 6 13 DM2
D4 14 6 DM2
VC 7 13 1.774
VE 14 4 1.774
IP 7 4 0.000374
DSUB 4 7 DM2
.MODEL QM1 NPN(IS=8e-16 BF=66670)
.MODEL QM2 NPN(IS=8.009E-16 BF=200000)
.MODEL DM1 D(IS=4.276E-12)
.MODEL DM2 D(IS=8e-16)
.ENDS LT1008
*-----------------------------------------------------------------------------
* connections: non-inverting input
* | inverting input
* | | positive power supply
* | | | negative power supply
* | | | | output
* | | | | | compensation
* | | | | | / \
.subckt LM301A 1 2 3 4 5 6 7
*
c1 11 12 8.661E-12
dc 5 53 dx
de 54 5 dx
dlp 90 91 dx
dln 92 90 dx
dp 4 3 dx
egnd 99 0 poly(2),(3,0),(4,0) 0 .5 .5
fb 7 99 poly(5) vb vc ve vlp vln 0 21.22E6 -20E6 20E6 20E6 -20E6
ga 6 0 11 12 188.5E-6
gcm 0 6 10 99 5.961E-9
iee 10 4 dc 15.14E-6
hlim 90 0 vlim 1K
q1 11 2 13 qx
q2 12 1 14 qx
r2 6 9 100.0E3
rc1 3 11 5.305E3
rc2 3 12 5.305E3
re1 13 10 1.839E3
re2 14 10 1.839E3
ree 10 99 13.21E6
ro1 8 5 50
ro2 7 99 25
rp 3 4 15.11E3
vb 9 0 dc 0
vc 3 53 dc 1
ve 54 4 dc 1
vlim 7 8 dc 0
vlp 91 0 dc 25
vln 0 92 dc 25
.model dx D(Is=800.0E-18 Rs=1)
.model qx NPN(Is=800.0E-18 Bf=107.1)
.ends
XU1 0 N006 N003 N007 N004 N002 N001 LM301A
V1 0 N007 15
V2 N003 0 15
V3 N005 0 SINE(0 1 1k)
R1 N004 N006 1k
R2 N006 N005 1k
C1 0 0 30p
.control
tran 50u 100m
run
print v(N004)
.endc